`default_nettype none `timescale 1ns / 1ns

module hazard_detector #(
    parameter logic [8:0] XLEN = 9'd64
) (
    input clk,
    input resetn
);

endmodule
