module led_blink (
input clk,
output reg led
);

// We want to blink an led here

endmodule
