`default_nettype none `timescale 1ns / 1ns

module uart_loopback_tb ();

initial begin
  $finish;
end

endmodule;
