`default_nettype none `timescale 1ns / 1ns

module riscv (
    input clk,
    input reset
);
endmodule
